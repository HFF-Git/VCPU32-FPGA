module MuxTB(


);

// fix .... see ChatGPT discussion ....

initial begin
    $dumpfile("@VCD_OUTPUT@");  // Placeholder for the VCD file name
    $dumpvars(0, your_top_module);
    // Other initialization code...
end



endmodule