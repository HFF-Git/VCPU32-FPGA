//------------------------------------------------------------------------------------------------------------
//
//  VCPU-32
//
//  Copyright (C) 2022 - 2024 Helmut Fieres, see License file.
//------------------------------------------------------------------------------------------------------------
// 
// - contains a lot of modules in one file...
// - test benches are however separate...
//
//
//------------------------------------------------------------------------------------------------------------
`ifndef PARAMETERS_VH
`define PARAMETERS_VH

// Common parameters for multiple modules
parameter int WIDTH = 8;
parameter int DEPTH = 256;
parameter int TIMEOUT = 100;

`endif // PARAMETERS_VH
