module MuxTB(


);

endmodule