module vcpu32(

    input logic clk
);

    always @( posedge clk ) begin

    end

endmodule


