//------------------------------------------------------------------------------------------------------------
//
//  VCPU-32
//
//  Copyright (C) 2022 - 2024 Helmut Fieres, see License file.
//------------------------------------------------------------------------------------------------------------
// 
// - contains a lot of modules in one file...
// - test benches are however separate...
//
//
//------------------------------------------------------------------------------------------------------------



//------------------------------------------------------------------------------------------------------------
//
//
//------------------------------------------------------------------------------------------------------------
`include "defines.vh"



//------------------------------------------------------------------------------------------------------------
//
//
//------------------------------------------------------------------------------------------------------------
module vcpu32(

    input logic clk
);

    register_file_16_32_3_2 U1 ( ); // example ....

    always @( posedge clk ) begin

    end

endmodule


