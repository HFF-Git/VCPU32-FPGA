//------------------------------------------------------------------------------------------------------------
//
//  VCPU-32
//
//  Copyright (C) 2022 - 2024 Helmut Fieres, see License file.
//------------------------------------------------------------------------------------------------------------
// 
// 
// - test benches are however separate...
//
//
//------------------------------------------------------------------------------------------------------------
`include "defines.vh"

//------------------------------------------------------------------------------------------------------------
//
//
//------------------------------------------------------------------------------------------------------------
module vcpu32(

    input logic     clk,
    input logic     rst

    );

    CpuCore CORE (  .clk( clk ), 
                    .rst( rst )
                        
                 );


    


    always @( negedge clk ) begin

    end

    always @( posedge clk ) begin

    end


endmodule


