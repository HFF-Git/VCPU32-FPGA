module vcpu32(


);



endmodule


